14 uid=262235
20 atime=1550777995
